pBAV       �o �� = / @  ���� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������  @$       �����  , � � � �   @%       �����  # � � � �   @&       �����   � � � �   @'       �����   � � � �   @(       �����   � � � �   @)       �����   � � � �   @*       �����   � � � �   @7       �����   � � � �   @,         �����  $ � � � �   @- !!      �����  % � � � �   @: ""      �����  & � � � �   @; ##      �����  ' � � � �   @< $$      �����  ( � � � �   @= %%      �����  ) � � � �   @> &&      �����  * � � � �   @? ''      �����  + � � � �   @$       ����� - � � � �   @%       ����� . � � � �   @&       �����   � � � �   @'       ����� ! � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       ����� / � � � �   @%       �����  � � � �   @&       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       ����� / � � � �   @%       �����  � � � �   @&       ����� 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       �����  � � � �   @%       �����  � � � �   @&       �����  � � � �   @'       �����  � � � �   @(       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       �����  � � � �   @%       �����  � � � �   @&       �����  � � � �   @'       �����  � � � �   @(       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       �����  � � � �   @%       �����  � � � �   @&       �����  � � � �   @'       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       �����  � � � �   @%       �����  � � � �   @&       �����  � � � �   @'       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       ����� 
 � � � �   @%       �����  � � � �   @&       �����  � � � �   @'       �����  � � � �   @(       �����  � � � �   @)       �����  � � � �   @*       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @$       �����	 
 � � � �   @%       �����	  � � � �   @&       �����	  � � � �   @'       �����	  � � � �   @(       �����	  � � � �   @)       �����	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �   @$       �����
  � � � �   @%       �����
  � � � �   @&       �����
  � � � �   @'       �����
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �      �|v(��z�������F��x��J�PF��;�h���br $ X r 6 �
$V                                                                                                                                                                                                                                                                                                                                                                                                                                